../Cap_voltage_v1_0/CapVoltage.vhd