../Profile_Sweep_v1_0/ProfileSweep.vhd