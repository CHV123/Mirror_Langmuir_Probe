../Div_int_delay_v1_0/DivIntDelay.vhd