../../../probe-response-current/cores/current_response_v1_0/CurRes.vhd