../current_response_v1_0/CurrentResponse.vhd