../Div_to_address_v1_0/DivToAdress.vhd