../input_control_v1_0/InputControl.vhd